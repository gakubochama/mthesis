module m_ALU();

endmodule

module m_decoder();

endmodule

module m_regfile();

endmodule

module m_shiftreg();

endmodule

module m_datapath();

endmodule